`include "modules/constants.v"

module notes_rom(
    input [1:0] noteType,
    input [4:0] addr,
    output reg [`NOTE_WIDTH-1:0] data
);
    always @(noteType, addr)
        case (noteType)
            `QUARTER_NOTE: case (addr)
                5'd00: data = 28'b0000000000000111111111110000;
                5'd01: data = 28'b0000000000011111111111111100;
                5'd02: data = 28'b0000000001111111111111111110;
                5'd03: data = 28'b0000000111111111111111111110;
                5'd04: data = 28'b0000001111111111111111111111;
                5'd05: data = 28'b0000011111111111111111111111;
                5'd06: data = 28'b0000111111111111111111111111;
                5'd07: data = 28'b0001111111111111111111111111;
                5'd08: data = 28'b0011111111111111111111111111;
                5'd09: data = 28'b0011111111111111111111111111;
                5'd10: data = 28'b0111111111111111111111111111;
                5'd11: data = 28'b0111111111111111111111111111;
                5'd12: data = 28'b1111111111111111111111111110;
                5'd13: data = 28'b1111111111111111111111111110;
                5'd14: data = 28'b1111111111111111111111111100;
                5'd15: data = 28'b1111111111111111111111111100;
                5'd16: data = 28'b1111111111111111111111111000;
                5'd17: data = 28'b1111111111111111111111110000;
                5'd18: data = 28'b1111111111111111111111100000;
                5'd19: data = 28'b1111111111111111111111000000;
                5'd20: data = 28'b0111111111111111111110000000;
                5'd21: data = 28'b0111111111111111111000000000;
                5'd22: data = 28'b0011111111111111100000000000;
                5'd23: data = 28'b0000111111111110000000000000;
            endcase
            `HALF_NOTE: case (addr)
                5'd00: data = 28'b0000000000000111111111110000;
                5'd01: data = 28'b0000000000011111111111111100;
                5'd02: data = 28'b0000000001111111111111111110;
                5'd03: data = 28'b0000000111111111111111111110;
                5'd04: data = 28'b0000001111111111111100001111;
                5'd05: data = 28'b0000011111111111100000000111;
                5'd06: data = 28'b0000111111111110000000000111;
                5'd07: data = 28'b0001111111111000000000001111;
                5'd08: data = 28'b0011111111110000000000001111;
                5'd09: data = 28'b0011111111000000000000011111;
                5'd10: data = 28'b0111111110000000000000111111;
                5'd11: data = 28'b0111111100000000000001111111;
                5'd12: data = 28'b1111111000000000000011111110;
                5'd13: data = 28'b1111110000000000000111111110;
                5'd14: data = 28'b1111100000000000001111111100;
                5'd15: data = 28'b1111000000000000111111111100;
                5'd16: data = 28'b1111000000000001111111111000;
                5'd17: data = 28'b1110000000000111111111110000;
                5'd18: data = 28'b1110000000011111111111100000;
                5'd19: data = 28'b1111000011111111111111000000;
                5'd20: data = 28'b0111111111111111111110000000;
                5'd21: data = 28'b0111111111111111111000000000;
                5'd22: data = 28'b0011111111111111100000000000;
                5'd23: data = 28'b0000111111111110000000000000;
            endcase
            `WHOLE_NOTE: case (addr)
                5'd00: data = 28'b0000000011111111111100000000;
                5'd01: data = 28'b0000001111111111111111000000;
                5'd02: data = 28'b0000111111111111111111110000;
                5'd03: data = 28'b0001111111000011111111111000;
                5'd04: data = 28'b0011111110000001111111111100;
                5'd05: data = 28'b0111111110000000111111111110;
                5'd06: data = 28'b0111111100000000011111111110;
                5'd07: data = 28'b1111111100000000011111111111;
                5'd08: data = 28'b1111111100000000001111111111;
                5'd09: data = 28'b1111111100000000001111111111;
                5'd10: data = 28'b1111111100000000000111111111;
                5'd11: data = 28'b1111111100000000000111111111;
                5'd12: data = 28'b1111111110000000000011111111;
                5'd13: data = 28'b1111111110000000000011111111;
                5'd14: data = 28'b1111111111000000000011111111;
                5'd15: data = 28'b1111111111000000000011111111;
                5'd16: data = 28'b1111111111100000000011111111;
                5'd17: data = 28'b0111111111100000000011111110;
                5'd18: data = 28'b0111111111110000000111111110;
                5'd19: data = 28'b0011111111111000000111111100;
                5'd20: data = 28'b0001111111111100001111111000;
                5'd21: data = 28'b0000111111111111111111110000;
                5'd22: data = 28'b0000001111111111111111000000;
                5'd23: data = 28'b0000000011111111111100000000;
            endcase
        endcase

endmodule
